library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;



entity nasobicka is
   Port ( 
      d : in  STD_LOGIC;
      c : in  STD_LOGIC; 
      b : in  STD_LOGIC;
      a : in  STD_LOGIC;
      outa : out  STD_LOGIC;
      outb : out  STD_LOGIC;
      outc : out  STD_LOGIC;
      outd : out  STD_LOGIC
   );
end nasobicka;                                       
-- popis chov�n� 7-segmentov�ho dekod�ru
architecture nasobicka_arch of nasobicka is       
   -- vnit�n� sign�l, kter� se pou��v� k rozli�en� jednotliv�ch vstup�
   signal   input :  std_logic_vector (3 downto 0);     
   
begin

   -- zpracov�n� vstup� pro jednodu��� pr�ci s tabulkou 
   input(3) <= d;
   input(2) <= c;
   input(1) <= b;
   input(0) <= a;
	

	
   -- ------------------------------------------------------------------------------
   -- |  fun�kn� hodnota cd(d, c, b, a) |  stavov� index s  |  d  |  c  |  b  |  a  | 
   -- ------------------------------------------------------------------------------
   with input select
   outd <= '0'   when	"0000",         -- |           0       |  0  |  0  |  0  |  0  |       
         '0'   when	"0001",         -- |           1       |  0  |  0  |  0  |  1  |
         '0'   when	"0010",         -- |           2       |  0  |  0  |  1  |  0  |
         '0'   when	"0011",         -- |           3       |  0  |  0  |  1  |  1  |
         '0'   when	"0100",         -- |           4       |  0  |  1  |  0  |  0  |
         '0'   when	"0101",         -- |           5       |  0  |  1  |  0  |  1  |
         '0'   when	"0110",         -- |           6       |  0  |  1  |  1  |  0  |
         '0'   when	"0111",         -- |           7       |  0  |  1  |  1  |  1  |
         '0'   when	"1000",         -- |           8       |  1  |  0  |  0  |  0  |
         '0'   when	"1001",         -- |           9       |  1  |  0  |  0  |  1  |
         '0'   when	"1010",         -- |          10 (A)   |  1  |  0  |  1  |  0  |
         '0'   when	"1011",         -- |          11 (b)   |  1  |  0  |  1  |  1  |
         '0'   when	"1100",         -- |          12 (C)   |  1  |  1  |  0  |  0  |
         '0'   when	"1101",         -- |          13 (d)   |  1  |  1  |  0  |  1  |
         '0'   when	"1110",         -- |          14 (E)   |  1  |  1  |  1  |  0  |
         '1'   when	"1111",         -- |          15 (F)   |  1  |  1  |  1  |  1  |
         '1'	when others;
   
   -- ------------------------------------------------------------------------------;
   -- ------------------------------------------------------------------------------
   -- |  fun�kn� hodnota ce(d, c, b, a) |  stavov� index s  |  d  |  c  |  b  |  a  | 
   -- ------------------------------------------------------------------------------
   with input select
   outc <= '0'   when	"0000",         -- |           0       |  0  |  0  |  0  |  0  |  
         '0'   when	"0001",         -- |           1       |  0  |  0  |  0  |  1  |   
         '0'   when	"0010",         -- |           2       |  0  |  0  |  1  |  0  |           
         '0'   when	"0011",         -- |           3       |  0  |  0  |  1  |  1  |
         '0'   when	"0100",         -- |           4       |  0  |  1  |  0  |  0  |   
         '0'   when	"0101",         -- |           5       |  0  |  1  |  0  |  1  |   
         '0'   when	"0110",         -- |           6       |  0  |  1  |  1  |  0  |
         '0'   when	"0111",         -- |           7       |  0  |  1  |  1  |  1  |
         '0'   when	"1000",         -- |           8       |  1  |  0  |  0  |  0  |
         '0'   when	"1001",         -- |           9       |  1  |  0  |  0  |  1  |
         '1'   when	"1010",         -- |          10 (A)   |  1  |  0  |  1  |  0  |
         '1'   when	"1011",         -- |          11 (b)   |  1  |  0  |  1  |  1  |
         '0'   when	"1100",         -- |          12 (C)   |  1  |  1  |  0  |  0  |
         '0'   when	"1101",         -- |          13 (d)   |  1  |  1  |  0  |  1  |
         '1'   when	"1110",         -- |          14 (E)   |  1  |  1  |  1  |  0  |
         '0'   when	"1111",         -- |          15 (F)   |  1  |  1  |  1  |  1  |
         '1'	when others;
   
   -- ------------------------------------------------------------------------------;
   -- ------------------------------------------------------------------------------
   -- |  fun�kn� hodnota cf(d, c, b, a) |  stavov� index s  |  d  |  c  |  b  |  a  | 
   -- ------------------------------------------------------------------------------
   with input select
   outb <= '0'   when	"0000",         -- |           0       |  0  |  0  |  0  |  0  |            
         '0'   when	"0001",         -- |           1       |  0  |  0  |  0  |  1  |
         '0'   when	"0010",         -- |           2       |  0  |  0  |  1  |  0  |
         '0'   when	"0011",         -- |           3       |  0  |  0  |  1  |  1  |
         '0'   when	"0100",         -- |           4       |  0  |  1  |  0  |  0  |           
         '0'   when	"0101",         -- |           5       |  0  |  1  |  0  |  1  |
         '1'   when	"0110",         -- |           6       |  0  |  1  |  1  |  0  |             
         '1'   when	"0111",         -- |           7       |  0  |  1  |  1  |  1  |           
         '0'   when	"1000",         -- |           8       |  1  |  0  |  0  |  0  |          
         '1'   when	"1001",         -- |           9       |  1  |  0  |  0  |  1  |          
         '0'   when	"1010",         -- |          10 (A)   |  1  |  0  |  1  |  0  |
         '1'   when	"1011",         -- |          11 (b)   |  1  |  0  |  1  |  1  |
         '0'   when	"1100",         -- |          12 (C)   |  1  |  1  |  0  |  0  |
         '1'   when	"1101",         -- |          13 (d)   |  1  |  1  |  0  |  1  |
         '1'   when	"1110",         -- |          14 (E)   |  1  |  1  |  1  |  0  |
         '0'   when	"1111",         -- |          15 (F)   |  1  |  1  |  1  |  1  |
         '1'	when others;
   
   -- ------------------------------------------------------------------------------;
   -- ------------------------------------------------------------------------------
   -- |  fun�kn� hodnota cg(d, c, b, a) |  stavov� index s  |  d  |  c  |  b  |  a  | 
   -- ------------------------------------------------------------------------------
   with input select
   outa <= '0'   when	"0000",         -- |           0       |  0  |  0  |  0  |  0  |     
         '0'   when	"0001",         -- |           1       |  0  |  0  |  0  |  1  |            
         '0'   when	"0010",         -- |           2       |  0  |  0  |  1  |  0  |         
         '0'   when	"0011",         -- |           3       |  0  |  0  |  1  |  1  |
         '0'   when	"0100",         -- |           4       |  0  |  1  |  0  |  0  |
         '1'   when	"0101",         -- |           5       |  0  |  1  |  0  |  1  |
         '0'   when	"0110",         -- |           6       |  0  |  1  |  1  |  0  |
         '1'   when	"0111",         -- |           7       |  0  |  1  |  1  |  1  |             
         '0'   when	"1000",         -- |           8       |  1  |  0  |  0  |  0  |             
         '0'   when	"1001",         -- |           9       |  1  |  0  |  0  |  1  |
         '0'   when	"1010",         -- |          10 (A)   |  1  |  0  |  1  |  0  |
         '0'   when	"1011",         -- |          11 (b)   |  1  |  0  |  1  |  1  |
         '0'   when	"1100",         -- |          12 (C)   |  1  |  1  |  0  |  0  |
         '1'   when	"1101",         -- |          13 (d)   |  1  |  1  |  0  |  1  |
         '0'   when	"1110",         -- |          14 (E)   |  1  |  1  |  1  |  0  |
         '1'   when	"1111",         -- |          15 (F)   |  1  |  1  |  1  |  1  |
         '1'	when others;
    
   -- ------------------------------------------------------------------------------;


	
end nasobicka_arch;

